module _and(
    input A,
    input B,
    output reg C
);

assign C = A & B;

endmodule