module add(
    input [3:0] A, B,
    output [3:0] Salida
);

assign Salida = A + B;

endmodule